`define PIPE
